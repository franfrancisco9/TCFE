* T3

* forces current values to be saved
.options savecurrents

Vin 3 1 DC 0 SIN(0  14.64891221288435 50 0 0 90)

*Envelop Detector

D1 0 3 default
D2 3 2 default
D3 1 2 default
D4 0 1 default

R1 2 0 26k

C 2 0 33.75u

*Voltage Regulator

R2 2 4 10k
Dr 4 0 Dmine
.MODEL Default D
.MODEL Dmine D (N=20)




* Transient simulation:
.control

set hcopypscolor=1
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=violet
set color5=rgb:3/8/0
set color6=rgb:4/0/0

op


tran 1e-5 0.2 0.0

plot  v(2)
hardcopy venv.eps v(2)


plot  v(4)
hardcopy vout.eps v(4)


plot v(4)-12
hardcopy vout(ac+dc).eps v(4)-12


plot v(1)-v(3) v(2) v(4)
hardcopy vs_vout.eps v(1)-v(3) v(2) 12 v(4) 

meas tran Output_average AVG v(4) 
meas tran Max MAX v(4)
meas tran Min MIN v(4) 

let ripple = Max - Min

print Output_average ripple

print 1/ (72.150* ((maximum(v(4))-minimum(v(4))) + abs(mean(v(4)-12)) + 10e-6))


quit
.endc
.end
