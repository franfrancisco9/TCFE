* T3

* forces current values to be saved
.options savecurrents

Vin 3 1 DC 0 SIN(0  230.1 50 0 0 90)

*Envelop Detector

D1 0 3 default
D2 3 2 default
D3 1 2 default
D4 0 1 default

R1 2 0 920k

C 2 0 920u

*Voltage Regulator

R2 2 4 30.3k
Dr 4 0 Dmine
.MODEL Default D
.MODEL Dmine D (N=17)




* Transient simulation:
.control

set hcopypscolor=1
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=violet
set color5=rgb:3/8/0
set color6=rgb:4/0/0

op


tran 1e-5 0.2 0.0

plot  v(2)
hardcopy venv.ps v(2)


plot  v(4)
hardcopy vout.ps v(4)


plot v(4)-12
hardcopy vout(ac+dc).ps v(4)-12


plot v(1)-v(3) v(2) v(4)
hardcopy vs_vout.ps v(1)-v(3) v(2) 12 v(4) 
echo vs_vout_FIG

meas tran Output_average AVG v(4) 
meas tran Max MAX v(4)
meas tran Min MIN v(4) 

let ripple = Max - Min

print Output_average ripple

print 1/ (1877.5* ((maximum(v(4))-minimum(v(4))) + abs(mean(v(4)-12)) + 10e-6))


quit
.endc
.end
