*voltage divider netlist
.options savecurrents

*.include ../mat/ngspice_circuit_1.txt
.include ../doc/ngspice_circuit_1.txt


.control

op

echo "********************************************"
echo  "Operating point"
echo "********************************************"

echo  "op_TAB"
print all
echo  "op_END"

echo "********************************************"
echo  "Given Values"
echo "********************************************"

echo "op_TAB1"
echo "R1 = 1.01949191994 KΩ" 
echo "R2 = 2.05054429461 KΩ"
echo "R3 = 3.09286027724 KΩ"
echo "R4 = 4.12838973576 KΩ"
echo "R5 = 3.06635427647 KΩ"
echo "R6 = 2.01254230153 KΩ"
echo "R7 = 1.00502981701 KΩ"
echo "Va = 5.24204797361 V"
echo "C = 1.01905568201 uF"
echo "Kb = 7.23185131759 mS"
echo "Kd = 8.12820254987 KΩ"
echo "op_END1"

quit

.endc 


*R1 = 1.01949191994 
*R2 = 2.05054429461 
*R3 = 3.09286027724 
*R4 = 4.12838973576 
*R5 = 3.06635427647 
*R6 = 2.01254230153 
*R7 = 1.00502981701 
*Vs = 5.24204797361 
*C = 1.01905568201 
*Kb = 7.23185131759 
*Kc = 8.12820254987

.end




