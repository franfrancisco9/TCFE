*-----------------------------------------------------------------------------
*
* To use a subcircuit, the name must begin with 'X'.  For example:
* X1 1 2 3 4 5 uA741
*
* connections:   non-inverting input
*                |  inverting input
*                |  |  positive power supply
*                |  |  |  negative power supply
*                |  |  |  |  output
*                |  |  |  |  |
.subckt uA741    1  2  3  4  5
*
  c1   11 12 8.661E-12
  c2    6  7 30.00E-12
  dc    5 53 dx
  de   54  5 dx
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2) (3,0) (4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 10.61E6 -10E6 10E6 10E6 -10E6
  ga    6  0 11 12 188.5E-6
  gcm   0  6 10 99 5.961E-9
  iee  10  4 dc 15.16E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 5.305E3
  rc2   3 12 5.305E3
  re1  13 10 1.836E3
  re2  14 10 1.836E3
  ree  10 99 13.19E6
  ro1   8  5 50
  ro2   7 99 100
  rp    3  4 18.16E3
  vb    9  0 dc 0
  vc    3 53 dc 1
  ve   54  4 dc 1
  vlim  7  8 dc 0
  vlp  91  0 dc 40
  vln   0 92 dc 40
.model dx D(Is=800.0E-18 Rs=1)
.model qx NPN(Is=800.0E-18 Bf=93.75)
.ends



.options savecurrents

Vcc vcc 0 10.0
Vee vee 0 -10.0
Vin vin 0 0 ac 1.0 sin(0 10m 1k)

X1 in_p inv_in vcc vee out uA741

* non-inv +
C1 vin in_p 220n
R1 in_p 0 1k

* inv -
R3 inv_in r3b 100k
R3b r3b out 100k
R3c r3b out 100k

R4 inv_in 0 1k

* load
R2 out vo 1k
C2 vo 0 110n

.op
.end

.control

*makes plots in color
set hcopypscolor=0
set color0=white
set color1=black
set color2=red
set color3=rgb:0/9/9
set color4=violet
set color5=rgb:3/8/0
set color6=rgb:4/0/0



*op
*print all

* time analysis
*tran 1e-5 1e-2
*plot v(out)
*hardcopy lab-vo1.ps v(vo) v(vin)
*print v(vin)[45] v(vo)[45]




echo ""
echo "**********************"
echo "* frequency analysis *"
echo "**********************"

ac dec 10 10 100MEG
*plot vdb(out)
*plot vp(out)
hardcopy lab-vo1f.ps vdb(vo) vp(vo)*180/pi


echo ""
echo "****************"
echo "* Cut-off Freq *"
echo "****************"

* cut-off freqs

let Av_db = vdb(vo)-vdb(vin)
meas ac voltGainDB MAX Av_db
let Av_m = vm(vo)/vm(vin)
meas ac voltGain MAX Av_m
let voltG3 = voltGainDB-3
*print voltG3

meas ac lowCOf WHEN Av_db=voltG3
meas ac Maxf MAX_AT Av_db
meas ac highCOf WHEN Av_db=voltG3 CROSS=LAST

let avgCOf = sqrt(lowCOf*highCOf)
print avgCOf

echo ""
echo "* op-amp *"
echo ""

let in_m = vm(in_p)/vm(vin)
meas ac inGain MAX in_m
let out_m = vm(out)/vm(vin)
meas ac outGain MAX out_m


echo ""
echo "*********"
echo "* merit *"
echo "*********"

let gain_deviation = abs(voltGainDB - 40)
let f_deviation = abs(avgCOf - 1k)
*let cost = 13323 + 
*let merit = 1/(cost*gain_deviation*f_deviation + 1/1000000)
print gain_deviation f_deviation 
*print cost merit

echo ""
echo "****************"
echo "* relative dev *"
echo "****************"

let gainperc = gain_deviation/40*100
let fperc = f_deviation/1k*100
print gainperc fperc


echo ""
echo "******************"
echo "* impedance ohm *"
echo "******************"
*input impedance in ohm
print abs(v(vin)[20]/vin#branch[20]/(-1))

let Zin = v(vin)[20]/vin#branch[20]/(-1)
let real=Re(Zin)
let imag=Im(Zin)
let absl=abs(Zin)


***************************** TABLES ******************************
echo ""
echo "**********"
echo "* TABLES *"
echo "**********"5 euros 

echo "inputZ_TAB"
echo "Zin = $&real + $&imag j"
echo " $|$\ Zin $|$\ = $&absl"
echo "inputZ_END"

let CentralFreq = avgCOf
let CentralFreqDev = f_deviation
let gainDeviation = gain_deviation
echo "merit_TAB"
print voltGainDB
print gainDeviation
print CentralFreq
print CentralFreqDev
*print cost
*print merit
print gainDeviation CentralFreqDev > results.txt
echo "merit_END"


echo "zin_TAB"
echo "$&absl"
echo "zin_END"

echo "gain1_TAB"
echo "$&voltGain"
echo "gain1_END"
echo "gain2_TAB"
echo "$&voltGainDB"
echo "gain2_END"

echo "freq1_TAB"
echo "$&lowCOf"
echo "freq1_END"
echo "freq2_TAB"
echo "$&highCOf"
echo "freq2_END"
echo "freq3_TAB"
echo "$&CentralFreq"
echo "freq3_END"

echo "percentages_TAB"
print gainperc fperc
echo "percentages_END"


*need a different setup to measure output impedance

quit
.endc 


