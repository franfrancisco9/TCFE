*voltage divider netlist
.options savecurrents

*.include ../mat/ngspice_circuit_2.txt
.include ../doc/ngspice_circuit_2.txt


.control

op

echo "********************************************"
echo  "Operating point 2"
echo "********************************************"

echo  "op_TAB2"
print all
echo  "op_END2"


quit

.endc 


*R1 = 1.01949191994 
*R2 = 2.05054429461 
*R3 = 3.09286027724 
*R4 = 4.12838973576 
*R5 = 3.06635427647 
*R6 = 2.01254230153 
*R7 = 1.00502981701 
*Vs = 5.24204797361 
*C = 1.01905568201 
*Kb = 7.23185131759 
*Kc = 8.12820254987

.end

