*voltage divider netlist
.options savecurrents

Va V1 V2 DC 5.24204797361 
R1 V6 V1 1.01949191994e+03
R2 V5 V6 2.05054429461e+03
R3 V6 V7 3.09286027724e+03
R4 V2 V7 4.12838973576e+03
R5 V4 V7 3.06635427647e+03
R6 V8 V3 2.01254230153e+03
R7 V3 0 1.00502981701e+03 
Id 0 V4 DC 1.01905568201e-03

*Vc
VVc V2 V8 0V
HVc V7 0 VVc 8.12820254987e+03 
*end Vc 

*Ib
GIb V4 V5 V6 V7 7.23185131759e-03
*end Ib

.control

op

echo "********************************************"
echo  "Operating point"
echo "********************************************"

echo  "op_TAB"
print all
echo  "op_END"

echo "********************************************"
echo  "Given Values"
echo "********************************************"

echo "op_TAB1"
echo "R1 = 1.01949191994 KΩ" 
echo "R2 = 2.05054429461 KΩ"
echo "R3 = 3.09286027724 KΩ"
echo "R4 = 4.12838973576 KΩ"
echo "R5 = 3.06635427647 KΩ"
echo "R6 = 2.01254230153 KΩ"
echo "R7 = 1.00502981701 KΩ"
echo "Va = 5.24204797361 V"
echo "Id = 1.01905568201 mA"
echo "Kb = 7.23185131759 mS"
echo "Kc = 8.12820254987 KΩ"
echo "op_END1"

quit 

.endc

*R1 = 1.01949191994 
*R2 = 2.05054429461 
*R3 = 3.09286027724 
*R4 = 4.12838973576 
*R5 = 3.06635427647 
*R6 = 2.01254230153 
*R7 = 1.00502981701 
*Vs = 5.24204797361 
*C = 1.01905568201 
*Kb = 7.23185131759 
*Kc = 8.12820254987

.end




