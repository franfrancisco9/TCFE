*Frequency response of Node 6
.options savecurrents

*.include ../mat/ngspice_circuit_5.txt
.include ../doc/ngspice_circuit_5.txt

.control

op


*makes plots in color
set hcopypscolor=0
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=violet
set color5=rgb:3/8/0
set color6=rgb:4/0/0

echo "********************************************"
echo  "Frequency analysis"
echo "********************************************"

ac dec 1000 0.1 1MEG



settype decibel out
hardcopy acm.eps vdb(V6) vdb(V1) xlimit 1 1000k ylabel 'small signal gain'
settype phase out

hardcopy acm1.eps cph(V6) cph(V1) xlimit 1 1000k ylabel 'phase (in rad)'

let outd(V6) = 180/PI*cph(V6) + 90
let outd(Vs) = 180/PI*cph(V1) + 90

settype phase outd
hardcopy acm2.eps outd(V6) outd(Vs) xlimit 1 1000k ylabel 'phase'



quit

.endc 


*R1 = 1.01949191994 
*R2 = 2.05054429461 
*R3 = 3.09286027724 
*R4 = 4.12838973576 
*R5 = 3.06635427647 
*R6 = 2.01254230153 
*R7 = 1.00502981701 
*Vs = 5.24204797361 
*C = 1.01905568201 
*Kb = 7.23185131759 
*Kc = 8.12820254987

.end



