*voltage divider netlist
.options savecurrents

*.include ../mat/ngspice_circuit_3.txt
.include ../doc/ngspice_circuit_3.txt

.control

op


echo "********************************************"
echo  "Transient analysis"
echo "********************************************"
tran 1e-5 20e-3 uic

*makes plots in color
set hcopypscolor=0
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=violet
set color5=rgb:3/8/0
set color6=rgb:4/0/0

hardcopy trans3.eps v(V6) 


quit

.endc 


*R1 = 1.01949191994 
*R2 = 2.05054429461 
*R3 = 3.09286027724 
*R4 = 4.12838973576 
*R5 = 3.06635427647 
*R6 = 2.01254230153 
*R7 = 1.00502981701 
*Vs = 5.24204797361 
*C = 1.01905568201 
*Kb = 7.23185131759 
*Kc = 8.12820254987

.end



