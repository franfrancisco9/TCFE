*voltage divider netlist
.options savecurrents

Vs V1 0 DC 5.24204797361
R1 V2 V1 1.01949191994e+03
R2 V3 V2 2.05054429461e+03
R3 V2 V5 3.09286027724e+03
R4 0 V5 4.12838973576e+03
R5 V6 V5 3.06635427647e+03
R6 V9 V7 2.01254230153e+03
R7 V7 V8 1.00502981701e+03 
Vx V6 V8  DC 8.763665


*Vc
VVc 0 V9 0V
HVc V5 V8 VVc 8.12820254987e+03 
*end Vc 

*Ib
GIb V6 V3 V2 V5 7.23185131759e-03
*end Ib

.control

op

echo "********************************************"
echo  "Operating point"
echo "********************************************"

echo  "op_TAB"
print all
echo  "op_END"

echo "********************************************"
echo  "Given Values"
echo "********************************************"

echo "op_TAB1"
echo "R1 = 1.01949191994 KΩ" 
echo "R2 = 2.05054429461 KΩ"
echo "R3 = 3.09286027724 KΩ"
echo "R4 = 4.12838973576 KΩ"
echo "R5 = 3.06635427647 KΩ"
echo "R6 = 2.01254230153 KΩ"
echo "R7 = 1.00502981701 KΩ"
echo "Va = 5.24204797361 V"
echo "C = 1.01905568201 F"
echo "Kb = 7.23185131759 mS"
echo "Kc = 8.12820254987 KΩ"
echo "op_END1"


quit

.endc 


*R1 = 1.01949191994 
*R2 = 2.05054429461 
*R3 = 3.09286027724 
*R4 = 4.12838973576 
*R5 = 3.06635427647 
*R6 = 2.01254230153 
*R7 = 1.00502981701 
*Vs = 5.24204797361 
*C = 1.01905568201 
*Kb = 7.23185131759 
*Kc = 8.12820254987

.end



